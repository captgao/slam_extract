`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2018/05/02 22:33:21
// Design Name: 
// Module Name: desc_compute
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module desc_compute(
    input clk,
    input start,
    input maskIn,

    input [247:0] col1,
    input [247:0] col2,
    input [247:0] col3,
    input [247:0] col4,
    input [247:0] col5,
    input [247:0] col6,
    input [247:0] col7,
    input [247:0] col8,
    input [247:0] col9,
    input [247:0] col10,
    input [247:0] col11,
    input [247:0] col12,
    input [247:0] col13,
    input [247:0] col14,
    input [247:0] col15,
    input [247:0] col16,
    input [247:0] col17,
    input [247:0] col18,
    input [247:0] col19,
    input [247:0] col20,
    input [247:0] col21,
    input [247:0] col22,
    input [247:0] col23,
    input [247:0] col24,
    input [247:0] col25,
    input [247:0] col26,
    input [247:0] col27,
    input [247:0] col28,
    input [247:0] col29,
    input [247:0] col30,
    input [247:0] col31,

    output [255:0] desc,
    output val,
    output maskOut

    );

    wire [7:0] src[0:255];
    wire [7:0] dst[0:255];
    reg [255:0] descReg = 0;
    reg valReg;

    assign desc = descReg;
    assign val = valReg;

    assign src[0]   =   col15[128:120];
    assign src[1]   =   col14[128:120];
    assign src[2]   =   col13[128:120];
    assign src[3]   =   col12[128:120];
    assign src[4]   =   col10[128:120];
    assign src[5]   =   col8[128:120];
    assign src[6]   =   col5[128:120];
    assign src[7]   =   col2[128:120];
    assign src[8]   =   col15[128:120];
    assign src[9]   =   col14[128:120];
    assign src[10]  =   col13[120:112];
    assign src[11]  =   col12[120:112];
    assign src[12]  =   col10[120:112];
    assign src[13]  =   col8[112:104];
    assign src[14]  =   col5[112:104];
    assign src[15]  =   col2[104:96];
    assign src[16]  =   col15[128:120];
    assign src[17]  =   col14[120:112];
    assign src[18]  =   col13[120:112];
    assign src[19]  =   col12[112:104];
    assign src[20]  =   col10[112:104];
    assign src[21]  =   col9[104:96];
    assign src[22]  =   col6[96:88];
    assign src[23]  =   col3[88:80];
    assign src[24]  =   col15[120:112];
    assign src[25]  =   col14[120:112];
    assign src[26]  =   col14[112:104];
    assign src[27]  =   col13[112:104];
    assign src[28]  =   col11[104:96];
    assign src[29]  =   col9[96:88];
    assign src[30]  =   col7[80:72];
    assign src[31]  =   col4[64:56];
    assign src[32]  =   col15[120:112];
    assign src[33]  =   col15[120:112];
    assign src[34]  =   col14[112:104];
    assign src[35]  =   col13[104:96];
    assign src[36]  =   col12[96:88];
    assign src[37]  =   col10[80:72];
    assign src[38]  =   col8[64:56];
    assign src[39]  =   col6[48:40];
    assign src[40]  =   col15[120:112];
    assign src[41]  =   col15[112:104];
    assign src[42]  =   col14[112:104];
    assign src[43]  =   col14[104:96];
    assign src[44]  =   col13[88:80];
    assign src[45]  =   col12[72:64];
    assign src[46]  =   col10[56:48];
    assign src[47]  =   col8[32:24];
    assign src[48]  =   col16[120:112];
    assign src[49]  =   col15[112:104];
    assign src[50]  =   col15[104:96];
    assign src[51]  =   col14[96:88];
    assign src[52]  =   col14[80:72];
    assign src[53]  =   col13[72:64];
    assign src[54]  =   col12[48:40];
    assign src[55]  =   col11[24:16];
    assign src[56]  =   col16[120:112];
    assign src[57]  =   col16[112:104];
    assign src[58]  =   col15[104:96];
    assign src[59]  =   col15[96:88];
    assign src[60]  =   col15[80:72];
    assign src[61]  =   col14[64:56];
    assign src[62]  =   col14[40:32];
    assign src[63]  =   col13[16:8];
    assign src[64]  =   col16[120:112];
    assign src[65]  =   col16[112:104];
    assign src[66]  =   col16[104:96];
    assign src[67]  =   col16[96:88];
    assign src[68]  =   col16[80:72];
    assign src[69]  =   col16[64:56];
    assign src[70]  =   col16[40:32];
    assign src[71]  =   col16[16:8];
    assign src[72]  =   col16[120:112];
    assign src[73]  =   col16[112:104];
    assign src[74]  =   col17[104:96];
    assign src[75]  =   col17[96:88];
    assign src[76]  =   col17[80:72];
    assign src[77]  =   col18[64:56];
    assign src[78]  =   col18[40:32];
    assign src[79]  =   col19[16:8];
    assign src[80]  =   col16[120:112];
    assign src[81]  =   col17[112:104];
    assign src[82]  =   col17[104:96];
    assign src[83]  =   col18[96:88];
    assign src[84]  =   col18[80:72];
    assign src[85]  =   col19[72:64];
    assign src[86]  =   col20[48:40];
    assign src[87]  =   col21[24:16];
    assign src[88]  =   col17[120:112];
    assign src[89]  =   col17[112:104];
    assign src[90]  =   col18[112:104];
    assign src[91]  =   col18[104:96];
    assign src[92]  =   col19[88:80];
    assign src[93]  =   col20[72:64];
    assign src[94]  =   col22[56:48];
    assign src[95]  =   col24[32:24];
    assign src[96]  =   col17[120:112];
    assign src[97]  =   col17[120:112];
    assign src[98]  =   col18[112:104];
    assign src[99]  =   col19[104:96];
    assign src[100] =   col20[96:88];
    assign src[101] =   col22[80:72];
    assign src[102] =   col24[64:56];
    assign src[103] =   col26[48:40];
    assign src[104] =   col17[120:112];
    assign src[105] =   col18[120:112];
    assign src[106] =   col18[112:104];
    assign src[107] =   col19[112:104];
    assign src[108] =   col21[104:96];
    assign src[109] =   col23[96:88];
    assign src[110] =   col25[80:72];
    assign src[111] =   col28[64:56];
    assign src[112] =   col17[128:120];
    assign src[113] =   col18[120:112];
    assign src[114] =   col19[120:112];
    assign src[115] =   col20[112:104];
    assign src[116] =   col22[112:104];
    assign src[117] =   col23[104:96];
    assign src[118] =   col26[96:88];
    assign src[119] =   col29[88:80];
    assign src[120] =   col17[128:120];
    assign src[121] =   col18[128:120];
    assign src[122] =   col19[120:112];
    assign src[123] =   col20[120:112];
    assign src[124] =   col22[120:112];
    assign src[125] =   col24[112:104];
    assign src[126] =   col27[112:104];
    assign src[127] =   col30[104:96];
    assign src[128] =   col17[128:120];
    assign src[129] =   col18[128:120];
    assign src[130] =   col19[128:120];
    assign src[131] =   col20[128:120];
    assign src[132] =   col22[128:120];
    assign src[133] =   col24[128:120];
    assign src[134] =   col27[128:120];
    assign src[135] =   col30[128:120];
    assign src[136] =   col17[128:120];
    assign src[137] =   col18[128:120];
    assign src[138] =   col19[136:128];
    assign src[139] =   col20[136:128];
    assign src[140] =   col22[136:128];
    assign src[141] =   col24[144:136];
    assign src[142] =   col27[144:136];
    assign src[143] =   col30[152:144];
    assign src[144] =   col17[128:120];
    assign src[145] =   col18[136:128];
    assign src[146] =   col19[136:128];
    assign src[147] =   col20[144:136];
    assign src[148] =   col22[144:136];
    assign src[149] =   col23[152:144];
    assign src[150] =   col26[160:152];
    assign src[151] =   col29[168:160];
    assign src[152] =   col17[136:128];
    assign src[153] =   col18[136:128];
    assign src[154] =   col18[144:136];
    assign src[155] =   col19[144:136];
    assign src[156] =   col21[152:144];
    assign src[157] =   col23[160:152];
    assign src[158] =   col25[176:168];
    assign src[159] =   col28[192:184];
    assign src[160] =   col17[136:128];
    assign src[161] =   col17[136:128];
    assign src[162] =   col18[144:136];
    assign src[163] =   col19[152:144];
    assign src[164] =   col20[160:152];
    assign src[165] =   col22[176:168];
    assign src[166] =   col24[192:184];
    assign src[167] =   col26[208:200];
    assign src[168] =   col17[136:128];
    assign src[169] =   col17[144:136];
    assign src[170] =   col18[144:136];
    assign src[171] =   col18[152:144];
    assign src[172] =   col19[168:160];
    assign src[173] =   col20[184:176];
    assign src[174] =   col22[200:192];
    assign src[175] =   col24[224:216];
    assign src[176] =   col16[136:128];
    assign src[177] =   col17[144:136];
    assign src[178] =   col17[152:144];
    assign src[179] =   col18[160:152];
    assign src[180] =   col18[176:168];
    assign src[181] =   col19[184:176];
    assign src[182] =   col20[208:200];
    assign src[183] =   col21[232:224];
    assign src[184] =   col16[136:128];
    assign src[185] =   col16[144:136];
    assign src[186] =   col17[152:144];
    assign src[187] =   col17[160:152];
    assign src[188] =   col17[176:168];
    assign src[189] =   col18[192:184];
    assign src[190] =   col18[216:208];
    assign src[191] =   col19[240:232];
    assign src[192] =   col16[136:128];
    assign src[193] =   col16[144:136];
    assign src[194] =   col16[152:144];
    assign src[195] =   col16[160:152];
    assign src[196] =   col16[176:168];
    assign src[197] =   col16[192:184];
    assign src[198] =   col16[216:208];
    assign src[199] =   col16[240:232];
    assign src[200] =   col16[136:128];
    assign src[201] =   col16[144:136];
    assign src[202] =   col15[152:144];
    assign src[203] =   col15[160:152];
    assign src[204] =   col15[176:168];
    assign src[205] =   col14[192:184];
    assign src[206] =   col14[216:208];
    assign src[207] =   col13[240:232];
    assign src[208] =   col16[136:128];
    assign src[209] =   col15[144:136];
    assign src[210] =   col15[152:144];
    assign src[211] =   col14[160:152];
    assign src[212] =   col14[176:168];
    assign src[213] =   col13[184:176];
    assign src[214] =   col12[208:200];
    assign src[215] =   col11[232:224];
    assign src[216] =   col15[136:128];
    assign src[217] =   col15[144:136];
    assign src[218] =   col14[144:136];
    assign src[219] =   col14[152:144];
    assign src[220] =   col13[168:160];
    assign src[221] =   col12[184:176];
    assign src[222] =   col10[200:192];
    assign src[223] =   col8[224:216];
    assign src[224] =   col15[136:128];
    assign src[225] =   col15[136:128];
    assign src[226] =   col14[144:136];
    assign src[227] =   col13[152:144];
    assign src[228] =   col12[160:152];
    assign src[229] =   col10[176:168];
    assign src[230] =   col8[192:184];
    assign src[231] =   col6[208:200];
    assign src[232] =   col15[136:128];
    assign src[233] =   col14[136:128];
    assign src[234] =   col14[144:136];
    assign src[235] =   col13[144:136];
    assign src[236] =   col11[152:144];
    assign src[237] =   col9[160:152];
    assign src[238] =   col7[176:168];
    assign src[239] =   col4[192:184];
    assign src[240] =   col15[128:120];
    assign src[241] =   col14[136:128];
    assign src[242] =   col13[136:128];
    assign src[243] =   col12[144:136];
    assign src[244] =   col10[144:136];
    assign src[245] =   col9[152:144];
    assign src[246] =   col6[160:152];
    assign src[247] =   col3[168:160];
    assign src[248] =   col15[128:120];
    assign src[249] =   col14[128:120];
    assign src[250] =   col13[136:128];
    assign src[251] =   col12[136:128];
    assign src[252] =   col10[136:128];
    assign src[253] =   col8[144:136];
    assign src[254] =   col5[144:136];
    assign src[255] =   col2[152:144];


    assign dst[0]   =   col21[128:120];
    assign dst[1]   =   col25[128:120];
    assign dst[2]   =   col20[128:120];
    assign dst[3]   =   col23[128:120];
    assign dst[4]   =   col29[128:120];
    assign dst[5]   =   col26[128:120];
    assign dst[6]   =   col19[128:120];
    assign dst[7]   =   col18[128:120];
    assign dst[8]   =   col21[136:128];
    assign dst[9]   =   col25[144:136];
    assign dst[10]  =   col20[136:128];
    assign dst[11]  =   col23[136:128];
    assign dst[12]  =   col29[152:144];
    assign dst[13]  =   col26[144:136];
    assign dst[14]  =   col19[136:128];
    assign dst[15]  =   col18[128:120];
    assign dst[16]  =   col21[144:136];
    assign dst[17]  =   col24[152:144];
    assign dst[18]  =   col20[144:136];
    assign dst[19]  =   col22[152:144];
    assign dst[20]  =   col28[168:160];
    assign dst[21]  =   col25[160:152];
    assign dst[22]  =   col19[136:128];
    assign dst[23]  =   col18[136:128];
    assign dst[24]  =   col20[152:144];
    assign dst[25]  =   col23[168:160];
    assign dst[26]  =   col19[144:136];
    assign dst[27]  =   col22[160:152];
    assign dst[28]  =   col27[184:176];
    assign dst[29]  =   col24[176:168];
    assign dst[30]  =   col18[144:136];
    assign dst[31]  =   col18[136:128];
    assign dst[32]  =   col20[160:152];
    assign dst[33]  =   col22[176:168];
    assign dst[34]  =   col19[152:144];
    assign dst[35]  =   col21[168:160];
    assign dst[36]  =   col25[200:192];
    assign dst[37]  =   col23[184:176];
    assign dst[38]  =   col18[144:136];
    assign dst[39]  =   col17[136:128];
    assign dst[40]  =   col19[160:152];
    assign dst[41]  =   col21[184:176];
    assign dst[42]  =   col18[152:144];
    assign dst[43]  =   col20[176:168];
    assign dst[44]  =   col23[216:208];
    assign dst[45]  =   col22[192:184];
    assign dst[46]  =   col18[144:136];
    assign dst[47]  =   col17[144:136];
    assign dst[48]  =   col18[168:160];
    assign dst[49]  =   col19[192:184];
    assign dst[50]  =   col18[160:152];
    assign dst[51]  =   col19[176:168];
    assign dst[52]  =   col21[224:216];
    assign dst[53]  =   col20[200:192];
    assign dst[54]  =   col17[152:144];
    assign dst[55]  =   col17[144:136];
    assign dst[56]  =   col17[168:160];
    assign dst[57]  =   col18[200:192];
    assign dst[58]  =   col17[160:152];
    assign dst[59]  =   col17[184:176];
    assign dst[60]  =   col19[232:224];
    assign dst[61]  =   col18[208:200];
    assign dst[62]  =   col17[152:144];
    assign dst[63]  =   col16[144:136];
    assign dst[64]  =   col16[168:160];
    assign dst[65]  =   col16[200:192];
    assign dst[66]  =   col16[160:152];
    assign dst[67]  =   col16[184:176];
    assign dst[68]  =   col16[232:224];
    assign dst[69]  =   col16[208:200];
    assign dst[70]  =   col16[152:144];
    assign dst[71]  =   col16[144:136];
    assign dst[72]  =   col15[168:160];
    assign dst[73]  =   col14[200:192];
    assign dst[74]  =   col15[160:152];
    assign dst[75]  =   col15[184:176];
    assign dst[76]  =   col13[232:224];
    assign dst[77]  =   col14[208:200];
    assign dst[78]  =   col15[152:144];
    assign dst[79]  =   col16[144:136];
    assign dst[80]  =   col14[168:160];
    assign dst[81]  =   col13[192:184];
    assign dst[82]  =   col14[160:152];
    assign dst[83]  =   col13[176:168];
    assign dst[84]  =   col11[224:216];
    assign dst[85]  =   col12[200:192];
    assign dst[86]  =   col15[152:144];
    assign dst[87]  =   col15[144:136];
    assign dst[88]  =   col13[160:152];
    assign dst[89]  =   col11[184:176];
    assign dst[90]  =   col14[152:144];
    assign dst[91]  =   col12[176:168];
    assign dst[92]  =   col9[216:208];
    assign dst[93]  =   col10[192:184];
    assign dst[94]  =   col14[144:136];
    assign dst[95]  =   col15[144:136];
    assign dst[96]  =   col12[160:152];
    assign dst[97]  =   col10[176:168];
    assign dst[98]  =   col13[152:144];
    assign dst[99]  =   col11[168:160];
    assign dst[100] =   col7[200:192];
    assign dst[101] =   col9[184:176];
    assign dst[102] =   col14[144:136];
    assign dst[103] =   col15[136:128];
    assign dst[104] =   col12[152:144];
    assign dst[105] =   col9[168:160];
    assign dst[106] =   col13[144:136];
    assign dst[107] =   col10[160:152];
    assign dst[108] =   col5[184:176];
    assign dst[109] =   col8[176:168];
    assign dst[110] =   col14[144:136];
    assign dst[111] =   col14[136:128];
    assign dst[112] =   col11[144:136];
    assign dst[113] =   col8[152:144];
    assign dst[114] =   col12[144:136];
    assign dst[115] =   col10[152:144];
    assign dst[116] =   col4[168:160];
    assign dst[117] =   col7[160:152];
    assign dst[118] =   col13[136:128];
    assign dst[119] =   col14[136:128];
    assign dst[120] =   col11[136:128];
    assign dst[121] =   col7[144:136];
    assign dst[122] =   col12[136:128];
    assign dst[123] =   col9[136:128];
    assign dst[124] =   col3[152:144];
    assign dst[125] =   col6[144:136];
    assign dst[126] =   col13[136:128];
    assign dst[127] =   col14[128:120];
    assign dst[128] =   col11[128:120];
    assign dst[129] =   col7[128:120];
    assign dst[130] =   col12[128:120];
    assign dst[131] =   col9[128:120];
    assign dst[132] =   col3[128:120];
    assign dst[133] =   col6[128:120];
    assign dst[134] =   col13[128:120];
    assign dst[135] =   col14[128:120];
    assign dst[136] =   col11[120:112];
    assign dst[137] =   col7[112:104];
    assign dst[138] =   col12[120:112];
    assign dst[139] =   col9[120:112];
    assign dst[140] =   col3[104:96];
    assign dst[141] =   col6[112:104];
    assign dst[142] =   col13[120:112];
    assign dst[143] =   col14[128:120];
    assign dst[144] =   col11[112:104];
    assign dst[145] =   col8[104:96];
    assign dst[146] =   col12[112:104];
    assign dst[147] =   col10[104:96];
    assign dst[148] =   col4[88:80];
    assign dst[149] =   col7[96:88];
    assign dst[150] =   col13[120:112];
    assign dst[151] =   col14[120:112];
    assign dst[152] =   col12[104:96];
    assign dst[153] =   col9[88:80];
    assign dst[154] =   col13[112:104];
    assign dst[155] =   col10[96:88];
    assign dst[156] =   col5[72:64];
    assign dst[157] =   col8[80:72];
    assign dst[158] =   col14[112:104];
    assign dst[159] =   col14[120:112];
    assign dst[160] =   col12[96:88];
    assign dst[161] =   col10[80:72];
    assign dst[162] =   col13[104:96];
    assign dst[163] =   col11[88:80];
    assign dst[164] =   col7[56:48];
    assign dst[165] =   col9[72:64];
    assign dst[166] =   col14[112:104];
    assign dst[167] =   col15[120:112];
    assign dst[168] =   col13[96:88];
    assign dst[169] =   col11[72:64];
    assign dst[170] =   col14[104:96];
    assign dst[171] =   col12[80:72];
    assign dst[172] =   col9[40:32];
    assign dst[173] =   col10[64:56];
    assign dst[174] =   col14[112:104];
    assign dst[175] =   col15[112:104];
    assign dst[176] =   col14[88:80];
    assign dst[177] =   col13[64:56];
    assign dst[178] =   col14[96:88];
    assign dst[179] =   col13[80:72];
    assign dst[180] =   col11[32:24];
    assign dst[181] =   col12[56:48];
    assign dst[182] =   col15[104:96];
    assign dst[183] =   col15[112:104];
    assign dst[184] =   col15[88:80];
    assign dst[185] =   col14[56:48];
    assign dst[186] =   col15[96:88];
    assign dst[187] =   col15[72:64];
    assign dst[188] =   col13[24:16];
    assign dst[189] =   col14[48:40];
    assign dst[190] =   col15[104:96];
    assign dst[191] =   col16[112:104];
    assign dst[192] =   col16[88:80];
    assign dst[193] =   col16[56:48];
    assign dst[194] =   col16[96:88];
    assign dst[195] =   col16[72:64];
    assign dst[196] =   col16[24:16];
    assign dst[197] =   col16[48:40];
    assign dst[198] =   col16[104:96];
    assign dst[199] =   col16[112:104];
    assign dst[200] =   col17[88:80];
    assign dst[201] =   col18[56:48];
    assign dst[202] =   col17[96:88];
    assign dst[203] =   col17[72:64];
    assign dst[204] =   col19[24:16];
    assign dst[205] =   col18[48:40];
    assign dst[206] =   col17[104:96];
    assign dst[207] =   col16[112:104];
    assign dst[208] =   col18[88:80];
    assign dst[209] =   col19[64:56];
    assign dst[210] =   col18[96:88];
    assign dst[211] =   col19[80:72];
    assign dst[212] =   col21[32:24];
    assign dst[213] =   col20[56:48];
    assign dst[214] =   col17[104:96];
    assign dst[215] =   col17[112:104];
    assign dst[216] =   col19[96:88];
    assign dst[217] =   col21[72:64];
    assign dst[218] =   col18[104:96];
    assign dst[219] =   col20[80:72];
    assign dst[220] =   col23[40:32];
    assign dst[221] =   col22[64:56];
    assign dst[222] =   col18[112:104];
    assign dst[223] =   col17[112:104];
    assign dst[224] =   col20[96:88];
    assign dst[225] =   col22[80:72];
    assign dst[226] =   col19[104:96];
    assign dst[227] =   col21[88:80];
    assign dst[228] =   col25[56:48];
    assign dst[229] =   col23[72:64];
    assign dst[230] =   col18[112:104];
    assign dst[231] =   col17[120:112];
    assign dst[232] =   col20[104:96];
    assign dst[233] =   col23[88:80];
    assign dst[234] =   col19[112:104];
    assign dst[235] =   col22[96:88];
    assign dst[236] =   col27[72:64];
    assign dst[237] =   col24[80:72];
    assign dst[238] =   col18[112:104];
    assign dst[239] =   col18[120:112];
    assign dst[240] =   col21[112:104];
    assign dst[241] =   col24[104:96];
    assign dst[242] =   col20[112:104];
    assign dst[243] =   col22[104:96];
    assign dst[244] =   col28[88:80];
    assign dst[245] =   col25[96:88];
    assign dst[246] =   col19[120:112];
    assign dst[247] =   col18[120:112];
    assign dst[248] =   col21[120:112];
    assign dst[249] =   col25[112:104];
    assign dst[250] =   col20[120:112];
    assign dst[251] =   col23[120:112];
    assign dst[252] =   col29[104:96];
    assign dst[253] =   col26[112:104];
    assign dst[254] =   col19[120:112];
    assign dst[255] =   col18[128:120];


    always@(posedge clk)
    begin
        valReg <= start;

        descReg[0] <= src[0]>dst[0];
        descReg[1] <= src[1]>dst[1];
        descReg[2] <= src[2]>dst[2];
        descReg[3] <= src[3]>dst[3];
        descReg[4] <= src[4]>dst[4];
        descReg[5] <= src[5]>dst[5];
        descReg[6] <= src[6]>dst[6];
        descReg[7] <= src[7]>dst[7];
        descReg[8] <= src[8]>dst[8];
        descReg[9] <= src[9]>dst[9];
        descReg[10] <= src[10]>dst[10];
        descReg[11] <= src[11]>dst[11];
        descReg[12] <= src[12]>dst[12];
        descReg[13] <= src[13]>dst[13];
        descReg[14] <= src[14]>dst[14];
        descReg[15] <= src[15]>dst[15];
        descReg[16] <= src[16]>dst[16];
        descReg[17] <= src[17]>dst[17];
        descReg[18] <= src[18]>dst[18];
        descReg[19] <= src[19]>dst[19];
        descReg[20] <= src[20]>dst[20];
        descReg[21] <= src[21]>dst[21];
        descReg[22] <= src[22]>dst[22];
        descReg[23] <= src[23]>dst[23];
        descReg[24] <= src[24]>dst[24];
        descReg[25] <= src[25]>dst[25];
        descReg[26] <= src[26]>dst[26];
        descReg[27] <= src[27]>dst[27];
        descReg[28] <= src[28]>dst[28];
        descReg[29] <= src[29]>dst[29];
        descReg[30] <= src[30]>dst[30];
        descReg[31] <= src[31]>dst[31];
        descReg[32] <= src[32]>dst[32];
        descReg[33] <= src[33]>dst[33];
        descReg[34] <= src[34]>dst[34];
        descReg[35] <= src[35]>dst[35];
        descReg[36] <= src[36]>dst[36];
        descReg[37] <= src[37]>dst[37];
        descReg[38] <= src[38]>dst[38];
        descReg[39] <= src[39]>dst[39];
        descReg[40] <= src[40]>dst[40];
        descReg[41] <= src[41]>dst[41];
        descReg[42] <= src[42]>dst[42];
        descReg[43] <= src[43]>dst[43];
        descReg[44] <= src[44]>dst[44];
        descReg[45] <= src[45]>dst[45];
        descReg[46] <= src[46]>dst[46];
        descReg[47] <= src[47]>dst[47];
        descReg[48] <= src[48]>dst[48];
        descReg[49] <= src[49]>dst[49];
        descReg[50] <= src[50]>dst[50];
        descReg[51] <= src[51]>dst[51];
        descReg[52] <= src[52]>dst[52];
        descReg[53] <= src[53]>dst[53];
        descReg[54] <= src[54]>dst[54];
        descReg[55] <= src[55]>dst[55];
        descReg[56] <= src[56]>dst[56];
        descReg[57] <= src[57]>dst[57];
        descReg[58] <= src[58]>dst[58];
        descReg[59] <= src[59]>dst[59];
        descReg[60] <= src[60]>dst[60];
        descReg[61] <= src[61]>dst[61];
        descReg[62] <= src[62]>dst[62];
        descReg[63] <= src[63]>dst[63];
        descReg[64] <= src[64]>dst[64];
        descReg[65] <= src[65]>dst[65];
        descReg[66] <= src[66]>dst[66];
        descReg[67] <= src[67]>dst[67];
        descReg[68] <= src[68]>dst[68];
        descReg[69] <= src[69]>dst[69];
        descReg[70] <= src[70]>dst[70];
        descReg[71] <= src[71]>dst[71];
        descReg[72] <= src[72]>dst[72];
        descReg[73] <= src[73]>dst[73];
        descReg[74] <= src[74]>dst[74];
        descReg[75] <= src[75]>dst[75];
        descReg[76] <= src[76]>dst[76];
        descReg[77] <= src[77]>dst[77];
        descReg[78] <= src[78]>dst[78];
        descReg[79] <= src[79]>dst[79];
        descReg[80] <= src[80]>dst[80];
        descReg[81] <= src[81]>dst[81];
        descReg[82] <= src[82]>dst[82];
        descReg[83] <= src[83]>dst[83];
        descReg[84] <= src[84]>dst[84];
        descReg[85] <= src[85]>dst[85];
        descReg[86] <= src[86]>dst[86];
        descReg[87] <= src[87]>dst[87];
        descReg[88] <= src[88]>dst[88];
        descReg[89] <= src[89]>dst[89];
        descReg[90] <= src[90]>dst[90];
        descReg[91] <= src[91]>dst[91];
        descReg[92] <= src[92]>dst[92];
        descReg[93] <= src[93]>dst[93];
        descReg[94] <= src[94]>dst[94];
        descReg[95] <= src[95]>dst[95];
        descReg[96] <= src[96]>dst[96];
        descReg[97] <= src[97]>dst[97];
        descReg[98] <= src[98]>dst[98];
        descReg[99] <= src[99]>dst[99];
        descReg[100] <= src[100]>dst[100];
        descReg[101] <= src[101]>dst[101];
        descReg[102] <= src[102]>dst[102];
        descReg[103] <= src[103]>dst[103];
        descReg[104] <= src[104]>dst[104];
        descReg[105] <= src[105]>dst[105];
        descReg[106] <= src[106]>dst[106];
        descReg[107] <= src[107]>dst[107];
        descReg[108] <= src[108]>dst[108];
        descReg[109] <= src[109]>dst[109];
        descReg[110] <= src[110]>dst[110];
        descReg[111] <= src[111]>dst[111];
        descReg[112] <= src[112]>dst[112];
        descReg[113] <= src[113]>dst[113];
        descReg[114] <= src[114]>dst[114];
        descReg[115] <= src[115]>dst[115];
        descReg[116] <= src[116]>dst[116];
        descReg[117] <= src[117]>dst[117];
        descReg[118] <= src[118]>dst[118];
        descReg[119] <= src[119]>dst[119];
        descReg[120] <= src[120]>dst[120];
        descReg[121] <= src[121]>dst[121];
        descReg[122] <= src[122]>dst[122];
        descReg[123] <= src[123]>dst[123];
        descReg[124] <= src[124]>dst[124];
        descReg[125] <= src[125]>dst[125];
        descReg[126] <= src[126]>dst[126];
        descReg[127] <= src[127]>dst[127];
        descReg[128] <= src[128]>dst[128];
        descReg[129] <= src[129]>dst[129];
        descReg[130] <= src[130]>dst[130];
        descReg[131] <= src[131]>dst[131];
        descReg[132] <= src[132]>dst[132];
        descReg[133] <= src[133]>dst[133];
        descReg[134] <= src[134]>dst[134];
        descReg[135] <= src[135]>dst[135];
        descReg[136] <= src[136]>dst[136];
        descReg[137] <= src[137]>dst[137];
        descReg[138] <= src[138]>dst[138];
        descReg[139] <= src[139]>dst[139];
        descReg[140] <= src[140]>dst[140];
        descReg[141] <= src[141]>dst[141];
        descReg[142] <= src[142]>dst[142];
        descReg[143] <= src[143]>dst[143];
        descReg[144] <= src[144]>dst[144];
        descReg[145] <= src[145]>dst[145];
        descReg[146] <= src[146]>dst[146];
        descReg[147] <= src[147]>dst[147];
        descReg[148] <= src[148]>dst[148];
        descReg[149] <= src[149]>dst[149];
        descReg[150] <= src[150]>dst[150];
        descReg[151] <= src[151]>dst[151];
        descReg[152] <= src[152]>dst[152];
        descReg[153] <= src[153]>dst[153];
        descReg[154] <= src[154]>dst[154];
        descReg[155] <= src[155]>dst[155];
        descReg[156] <= src[156]>dst[156];
        descReg[157] <= src[157]>dst[157];
        descReg[158] <= src[158]>dst[158];
        descReg[159] <= src[159]>dst[159];
        descReg[160] <= src[160]>dst[160];
        descReg[161] <= src[161]>dst[161];
        descReg[162] <= src[162]>dst[162];
        descReg[163] <= src[163]>dst[163];
        descReg[164] <= src[164]>dst[164];
        descReg[165] <= src[165]>dst[165];
        descReg[166] <= src[166]>dst[166];
        descReg[167] <= src[167]>dst[167];
        descReg[168] <= src[168]>dst[168];
        descReg[169] <= src[169]>dst[169];
        descReg[170] <= src[170]>dst[170];
        descReg[171] <= src[171]>dst[171];
        descReg[172] <= src[172]>dst[172];
        descReg[173] <= src[173]>dst[173];
        descReg[174] <= src[174]>dst[174];
        descReg[175] <= src[175]>dst[175];
        descReg[176] <= src[176]>dst[176];
        descReg[177] <= src[177]>dst[177];
        descReg[178] <= src[178]>dst[178];
        descReg[179] <= src[179]>dst[179];
        descReg[180] <= src[180]>dst[180];
        descReg[181] <= src[181]>dst[181];
        descReg[182] <= src[182]>dst[182];
        descReg[183] <= src[183]>dst[183];
        descReg[184] <= src[184]>dst[184];
        descReg[185] <= src[185]>dst[185];
        descReg[186] <= src[186]>dst[186];
        descReg[187] <= src[187]>dst[187];
        descReg[188] <= src[188]>dst[188];
        descReg[189] <= src[189]>dst[189];
        descReg[190] <= src[190]>dst[190];
        descReg[191] <= src[191]>dst[191];
        descReg[192] <= src[192]>dst[192];
        descReg[193] <= src[193]>dst[193];
        descReg[194] <= src[194]>dst[194];
        descReg[195] <= src[195]>dst[195];
        descReg[196] <= src[196]>dst[196];
        descReg[197] <= src[197]>dst[197];
        descReg[198] <= src[198]>dst[198];
        descReg[199] <= src[199]>dst[199];
        descReg[200] <= src[200]>dst[200];
        descReg[201] <= src[201]>dst[201];
        descReg[202] <= src[202]>dst[202];
        descReg[203] <= src[203]>dst[203];
        descReg[204] <= src[204]>dst[204];
        descReg[205] <= src[205]>dst[205];
        descReg[206] <= src[206]>dst[206];
        descReg[207] <= src[207]>dst[207];
        descReg[208] <= src[208]>dst[208];
        descReg[209] <= src[209]>dst[209];
        descReg[210] <= src[210]>dst[210];
        descReg[211] <= src[211]>dst[211];
        descReg[212] <= src[212]>dst[212];
        descReg[213] <= src[213]>dst[213];
        descReg[214] <= src[214]>dst[214];
        descReg[215] <= src[215]>dst[215];
        descReg[216] <= src[216]>dst[216];
        descReg[217] <= src[217]>dst[217];
        descReg[218] <= src[218]>dst[218];
        descReg[219] <= src[219]>dst[219];
        descReg[220] <= src[220]>dst[220];
        descReg[221] <= src[221]>dst[221];
        descReg[222] <= src[222]>dst[222];
        descReg[223] <= src[223]>dst[223];
        descReg[224] <= src[224]>dst[224];
        descReg[225] <= src[225]>dst[225];
        descReg[226] <= src[226]>dst[226];
        descReg[227] <= src[227]>dst[227];
        descReg[228] <= src[228]>dst[228];
        descReg[229] <= src[229]>dst[229];
        descReg[230] <= src[230]>dst[230];
        descReg[231] <= src[231]>dst[231];
        descReg[232] <= src[232]>dst[232];
        descReg[233] <= src[233]>dst[233];
        descReg[234] <= src[234]>dst[234];
        descReg[235] <= src[235]>dst[235];
        descReg[236] <= src[236]>dst[236];
        descReg[237] <= src[237]>dst[237];
        descReg[238] <= src[238]>dst[238];
        descReg[239] <= src[239]>dst[239];
        descReg[240] <= src[240]>dst[240];
        descReg[241] <= src[241]>dst[241];
        descReg[242] <= src[242]>dst[242];
        descReg[243] <= src[243]>dst[243];
        descReg[244] <= src[244]>dst[244];
        descReg[245] <= src[245]>dst[245];
        descReg[246] <= src[246]>dst[246];
        descReg[247] <= src[247]>dst[247];
        descReg[248] <= src[248]>dst[248];
        descReg[249] <= src[249]>dst[249];
        descReg[250] <= src[250]>dst[250];
        descReg[251] <= src[251]>dst[251];
        descReg[252] <= src[252]>dst[252];
        descReg[253] <= src[253]>dst[253];
        descReg[254] <= src[254]>dst[254];
        descReg[255] <= src[255]>dst[255];
    end

    reg maskReg = 0;
    always @(posedge clk)
        maskReg <= maskIn;
    
    assign maskOut = maskReg;

endmodule
